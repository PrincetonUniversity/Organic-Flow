VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "_<>" ;
DIVIDERCHAR "/" ;

MACRO NAND2X1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN NAND2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9250 BY 4100 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 8205 500 9150 995 ;
    END
    PORT
      LAYER M1 ;
        RECT 8105 400 9250 1095 ;
    END
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 4105 2555 5095 3545 ;
    END
    PORT
      LAYER M1 ;
        RECT 4105 2555 5095 3545 ;
    END
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7750 1300 8750 2000 ;
        RECT 7750 2300 8750 2860 ;
        RECT 5650 2300 6650 2860 ;
        RECT 5650 2000 8750 2300 ;
        RECT 5800 1440 5900 2000 ;
    END
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 4000 9250 4100 ;
    END
  END VDD

  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 0 0 9250 100 ;
    END
  END GND

  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 1250 9250 1350 ;
    END
  END VSS

  OBS
    LAYER M1 ;
      RECT 500 2300 1500 2860 ;
      RECT 500 2000 4600 2300 ;
      RECT 2600 2300 3600 2860 ;
      RECT 4100 1110 4600 2000 ;
      RECT 3250 1440 3350 2000 ;
      RECT 1500 500 3350 850 ;
        RECT 1505 850 2495 1695 ;
        RECT 3250 850 3350 1360 ;
        RECT 500 2940 1500 4100 ;
        RECT 2600 2940 3600 4100 ;
        RECT 5650 2940 6650 4100 ;
        RECT 7750 2940 8750 4100 ;
        RECT 5350 0 6350 100 ;
        RECT 5800 100 5900 1360 ;
    LAYER GA ;
      RECT 4100 1110 6850 1690 ;
      RECT 1500 1690 2500 1700 ;
      RECT 1500 1110 3850 1690 ;
      RECT 1500 700 2500 1110 ;
      RECT 7250 2610 9250 3190 ;
      RECT 9150 1000 9250 2610 ;
      RECT 8200 500 9250 1000 ;
      RECT 0 600 100 2610 ;
      RECT 0 2610 2000 3190 ;
      RECT 0 500 9250 600 ;
      RECT 2100 2610 7100 3190 ;
      RECT 4100 3190 5100 3550 ;
      RECT 4100 2550 5100 2610 ;
    LAYER CO ;
        RECT 1505 705 2495 1695 ;
      RECT 4105 1155 4595 1645 ;
    LAYER Via ;
        RECT 1800 1300 1810 1310 ;
        RECT 2000 1300 2010 1310 ;
        RECT 2200 1300 2210 1310 ;
        RECT 800 4050 810 4060 ;
        RECT 1000 4050 1010 4060 ;
        RECT 1200 4050 1210 4060 ;
        RECT 2900 4050 2910 4060 ;
        RECT 3100 4050 3110 4060 ;
        RECT 3300 4050 3310 4060 ;
        RECT 5900 4050 5910 4060 ;
        RECT 6100 4050 6110 4060 ;
        RECT 6300 4050 6310 4060 ;
        RECT 8000 4050 8010 4060 ;
        RECT 8300 4050 8310 4060 ;
        RECT 8500 4050 8510 4060 ;
        RECT 5650 45 5660 55 ;
        RECT 5850 45 5860 55 ;
        RECT 6050 45 6060 55 ;
  END
END NAND2X1

MACRO NOR2X1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN NOR2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9250 BY 4100 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 8205 500 9150 995 ;
    END
    PORT
      LAYER M1 ;
        RECT 8105 400 9250 1095 ;
    END
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 4105 2555 5095 3545 ;
    END
    PORT
      LAYER M1 ;
        RECT 4105 2555 5095 3545 ;
    END
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7750 1300 8750 2000 ;
        RECT 7750 2300 8750 2860 ;
        RECT 5650 2300 6650 2860 ;
        RECT 5650 2000 8750 2300 ;
        RECT 5800 1440 5900 2000 ;
    END
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 4000 9250 4100 ;
    END
  END VDD

  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 0 0 9250 100 ;
    END
  END GND

  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 1250 9250 1350 ;
    END
  END VSS

  OBS
    LAYER M1 ;
      RECT 500 2300 1500 2860 ;
      RECT 500 2000 4600 2300 ;
      RECT 2600 2300 3600 2860 ;
      RECT 4100 1110 4600 2000 ;
      RECT 3250 1440 3350 2000 ;
      RECT 1500 500 3350 850 ;
        RECT 1505 850 2495 1695 ;
        RECT 3250 850 3350 1360 ;
      RECT 500 2940 1500 4100 ;
        RECT 2600 2940 3600 4100 ;
        RECT 5650 2940 6650 4100 ;
        RECT 7750 2940 8750 4100 ;
        RECT 5350 0 6350 100 ;
        RECT 5800 100 5900 1360 ;
    LAYER GA ;
      RECT 4100 1110 6850 1690 ;
      RECT 1500 1690 2500 1700 ;
      RECT 1500 1110 3850 1690 ;
      RECT 1500 700 2500 1110 ;
      RECT 7250 2610 9250 3190 ;
      RECT 9150 1000 9250 2610 ;
      RECT 8200 500 9250 1000 ;
      RECT 0 600 100 2610 ;
      RECT 0 2610 2000 3190 ;
      RECT 0 500 9250 600 ;
      RECT 2100 2610 7100 3190 ;
      RECT 4100 3190 5100 3550 ;
      RECT 4100 2550 5100 2610 ;
    LAYER CO ;
      RECT 1505 705 2495 1695 ;
      RECT 4105 1155 4595 1645 ;
    LAYER Via ;
        RECT 1800 1300 1810 1310 ;
        RECT 2000 1300 2010 1310 ;
        RECT 2200 1300 2210 1310 ;
        RECT 800 4050 810 4060 ;
        RECT 1000 4050 1010 4060 ;
        RECT 1200 4050 1210 4060 ;
        RECT 2900 4050 2910 4060 ;
        RECT 3100 4050 3110 4060 ;
        RECT 3300 4050 3310 4060 ;
        RECT 5900 4050 5910 4060 ;
        RECT 6100 4050 6110 4060 ;
        RECT 6300 4050 6310 4060 ;
        RECT 8000 4050 8010 4060 ;
        RECT 8300 4050 8310 4060 ;
        RECT 8500 4050 8510 4060 ;
        RECT 5650 45 5660 55 ;
        RECT 5850 45 5860 55 ;
        RECT 6050 45 6060 55 ;

  END
END NOR2X1

MACRO INVX1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN INVX1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 5250 BY 4100 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 300 2870 1100 3670 ;
    END
    PORT
      LAYER M1 ;
        RECT 200 2770 1200 3770 ;
    END
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2950 1300 4050 1820 ;
        RECT 3650 1820 5200 2200 ;
        RECT 3650 2200 4650 2720 ;
    END
  END Y

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 4000 5200 4100 ;
    END
  END VDD

  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 0 0 5200 100 ;
    END
  END GND

  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 0 1250 5200 1350 ;
    END
  END VSS

  OBS
    LAYER M1 ;
      RECT 1735 1300 1835 1820 ;
      RECT 1735 1820 3000 2250 ;
      RECT 2700 1000 3000 1820 ;
      RECT 1800 2200 2800 2720 ;
      RECT 2700 1035 3290 1620 ;
      RECT 0 470 1000 1560 ;
      RECT 1000 470 1835 700 ;
      RECT 1735 700 1835 1200 ;
      RECT 1800 2820 2800 4100 ;
      RECT 3650 2820 4650 4100 ;
       RECT 3500 0 4500 100 ;
        RECT 3950 100 4050 1020 ;
    LAYER CO ;
        RECT 100 570 900 1460 ;
      RECT 2730 1135 3190 1520 ;
    LAYER Via ;
        RECT 300 1300 310 1310 ;
        RECT 500 1300 510 1310 ;
        RECT 800 1300 810 1310 ;
        RECT 2000 4050 2010 4060 ;
        RECT 2300 4050 2310 4060 ;
        RECT 2600 4050 2610 4060 ;
        RECT 3800 4050 3810 4060 ;
        RECT 4100 4050 4110 4060 ;
        RECT 4400 4050 4410 4060 ;
        RECT 3700 45 3710 55 ;
        RECT 4000 45 4010 55 ;
        RECT 4300 45 4310 55 ;
  END
END INVX1


END LIBRARY
