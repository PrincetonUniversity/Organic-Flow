.GLOBAL vdd vss vee 

.subckt __nand A B Y  length=10u w1=100u w2=20u w3=10u w4=10u
m1 4 A vdd vdd pmos l=length w=w1
m2 4 B vdd vdd pmos l=length w=w1
m3 Y A vdd vdd pmos l=length w=w2
m4 Y B vdd vdd pmos l=length w=w2
m5 vee vee 4 vdd pmos l=length w=w3
m6 vss 4 Y vdd pmos l=length w=w4
.ends __nand

.subckt NAND2X1 A B Y  
XI5 A B Y __nand 
.ends NAND2X1

