.GLOBAL vdd vss vee

.subckt __nand3 vout A B C length=10u w1=50u w2=30u w3=10u w4=10u
m1 4 A vdd vdd pmos l=length w=w1
m2 4 B vdd vdd pmos l=length w=w1
m3 4 C vdd vdd pmos l=length w=w1
m4 vout A vdd vdd pmos l=length w=w2
m5 vout B vdd vdd pmos l=length w=w2
m6 vout C vdd vdd pmos l=length w=w2
m7 vee vee 4 vdd pmos l=length w=w3
m8 vss 4 vout vdd pmos l=length w=w4
.ends __nand3

.subckt DFFASRX1 Q Qbar D CK PREbar CLRbar
X1 1 PREbar 4 2 __nand3
X2 2 1 CLRbar CK __nand3
X3 3 2 CK 4 __nand3
X4 4 3 CLRbar D __nand3
X5 Q PREbar 2 Qbar __nand3
X6 Qbar Q 3 CLRbar __nand3
.ends DFFASRX1